module top_module(zero);

    output zero;
    wire zero;
    assign zero=0;
    
endmodule